`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/13/2025 02:07:10 PM
// Design Name: 
// Module Name: Datapath
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Datapath( Clk);
   wire ReadRegister1, ReadRegister2, WriteRegister, WriteData, RegWrite, Clk, ReadData1,
    ReadData2, ALUControl, A, B, ALUResult, Zero,Address, WriteData, Clk, MemWrite, MemRead, ReadData,
    out, inA, inB, sel, in, out;
    
module RegisterFile(ReadRegister1, ReadRegister2, WriteRegister, WriteData, RegWrite, Clk, ReadData1, ReadData2);
module ALU32Bit(ALUControl, A, B, ALUResult, Zero);
module DataMemory(Address, WriteData, Clk, MemWrite, MemRead, ReadData); 
module Mux32Bit2To1(out, inA, inB, sel);
module SignExtension(in, out);
module Adder(AdderInput1,AdderInput2, AdderOutput );
module InstructionMemory(Address, Instruction); 

/////////////////////////F////////////////////////////////////////////////////////////////////////////////

/////////////////////////D//////////////////////////////////////////////////////////////////////////////

/////////////////////////E//////////////////////////////////////////////////////////////////////////////

/////////////////////////M//////////////////////////////////////////////////////////////////////////////

/////////////////////////W//////////////////////////////////////////////////////////////////////////////

endmodule
